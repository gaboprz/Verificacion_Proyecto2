//`timescale 1ns/1ps

// Incluir UVM
import uvm_pkg::*;
`include "uvm_macros.svh"

// Definiciones del proyecto
`include "mesh_defines.svh"

// Interfaces
`include "interface.sv"

// Componentes UVM
`include "sequence_item.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"

// DUT
`include "Router_library.sv"

module tb;

  // Señales globales
  logic clk;
  logic reset;

  // Señales para el DUT - arrays para `NUM_DEVS
  logic                      pndng[`NUM_DEVS];
  logic [`PKG_SZ-1:0]        data_out[`NUM_DEVS];
  logic                      popin[`NUM_DEVS];
  logic                      pop[`NUM_DEVS];
  logic [`PKG_SZ-1:0]        data_out_i_in[`NUM_DEVS];
  logic                      pndng_i_in[`NUM_DEVS];

  // Generación de reloj (100 MHz)
  initial begin
    clk = 1'b0;
    forever #5 clk = ~clk;  // período 10 ns
  end

  // Reset
  initial begin
    reset = 1'b1;
    #100 reset = 1'b0;
  end

  // Instanciación del DUT
  mesh_gnrtr #(
    .ROWS       (`ROWS),
    .COLUMS     (`COLUMNS),   // ← nombre del parámetro tal como está en el DUT
    .pckg_sz    (`PKG_SZ),
    .fifo_depth (`FIFO_DEPTH),
    .bdcst      (`BROADCAST)
  ) dut (
    .pndng        (pndng),
    .data_out     (data_out),
    .popin        (popin),
    .pop          (pop),
    .data_out_i_in(data_out_i_in),
    .pndng_i_in   (pndng_i_in),
    .clk          (clk),
    .reset        (reset)
  );

  // Interfaces virtuales para cada dispositivo
  router_external_if ext_if[`NUM_DEVS](clk, reset);

  // Conexión de interfaces al DUT
  generate
    for (genvar i = 0; i < `NUM_DEVS; i++) begin : connect_interfaces
      // TB -> DUT (entradas del DUT)
      assign data_out_i_in[i] = ext_if[i].data_out_i_in;
      assign pndng_i_in[i]    = ext_if[i].pndng_i_in;
      assign pop[i]           = ext_if[i].pop;

      // DUT -> TB (salidas del DUT)
      assign ext_if[i].data_out = data_out[i];
      assign ext_if[i].pndng    = pndng[i];
      assign ext_if[i].popin    = popin[i];
    end
  endgenerate

  // SINK simple para salida (el "consumidor" acepta cuando hay dato)
  generate
    for (genvar i = 0; i < `NUM_DEVS; i++) begin : auto_pop_sink
      always_ff @(posedge clk or posedge reset) begin
        if (reset) ext_if[i].pop <= 1'b0;
        else       ext_if[i].pop <= ext_if[i].pndng; // ready=1 cuando hay dato
      end
    end
  endgenerate

  // Registro de interfaces en config_db
  initial begin
    for (int i = 0; i < `NUM_DEVS; i++) begin
      string if_name = $sformatf("ext_if[%0d]", i);
      uvm_config_db#(virtual router_external_if)::set(null, "uvm_test_top.env.*", if_name, ext_if[i]);
      `uvm_info("TB", $sformatf("Interface %s registered", if_name), UVM_LOW)
    end
  end

  // Monitoreo básico del testbench
  initial begin
    #200; // Esperar a que termine el reset
    forever begin
      @(posedge clk);
      for (int i = 0; i < `NUM_DEVS; i++) begin
        if (pndng_i_in[i] === 1'b1) begin
          $display("[TB_MON] Time %0t: Device %0d sending packet: %h", 
                   $time, i, data_out_i_in[i]);
        end
        if (pndng[i] === 1'b1 && pop[i] === 1'b1) begin
          $display("[TB_MON] Time %0t: Device %0d received packet: %h", 
                   $time, i, data_out[i]);
        end
      end
    end
  end

  // Iniciar test UVM
  initial begin
    `uvm_info("TB", "Starting UVM test", UVM_LOW)
    run_test("base_test");
  end

  // Timeout
  initial begin
    #5000;  // 5 us
    `uvm_info("TB", "Timeout - finalizando simulación", UVM_LOW)
    $finish;
  end

  // Dump de waveforms (opcional)
  initial begin
    if ($test$plusargs("wave")) begin
      $dumpfile("mesh_waves.vcd");
      $dumpvars(0, tb);
      `uvm_info("TB", "Waveform dumping enabled", UVM_LOW)
    end
  end

endmodule