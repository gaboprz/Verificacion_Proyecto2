class gen_mesh_seq extends uvm_sequence;
  `uvm_object_utils(gen_mesh_seq)
  
  function new(string name="gen_mesh_seq");
    super.new(name);
  endfunction
  
  rand int num; 	// Número de paquetes a generar
  
  constraint c1 { num inside {[2:5]}; }
  
  virtual task body();
    for (int i = 0; i < num; i++) begin
      mesh_pkt m_item = mesh_pkt::type_id::create("m_item");
      start_item(m_item);
      m_item.randomize();
      `uvm_info("SEQ", $sformatf("Generate new item: %s", m_item.convert2str()), UVM_LOW)
      finish_item(m_item);
    end
    `uvm_info("SEQ", $sformatf("Done generation of %0d items", num), UVM_LOW)
  endtask
endclass