/////////////////////////////////////////////////////////////////////////////////////////////////////////
// Se define el sequence item
/////////////////////////////////////////////////////////////////////////////////////////////////////////

`include "mesh_defines.svh"

class mesh_pkt extends uvm_sequence_item;
  `uvm_object_utils(mesh_pkt)

  // Campos del paquete
  rand bit [7:0]            nxt_jump;
  rand bit [3:0]            target_row;
  rand bit [3:0]            target_col;
  rand bit                  mode;
  rand bit [`PAYLOAD_W-1:0] payload;

  // Vector listo para el DUT
  bit [`PKG_SZ-1:0]         raw_pkt;

  // (nuevo) puerto de salida observado por el monitor (no rand)
  int unsigned              egress_id;

  // Constraints
  constraint c_nxt_no_bcast { nxt_jump != 8'hFF; }
  constraint c_row { target_row inside {[0:`ROWS-1]}; }
  constraint c_col { target_col inside {[0:`COLUMNS-1]}; }

  function new(string name="mesh_pkt"); super.new(name); endfunction

  function void pack_bits();
    raw_pkt = '0;
    raw_pkt[`PKG_SZ-1   -: 8]  = nxt_jump;
    raw_pkt[`PKG_SZ-9   -: 4]  = target_row;
    raw_pkt[`PKG_SZ-13  -: 4]  = target_col;
    raw_pkt[`PKG_SZ-17]        = mode;
    if (`PAYLOAD_W > 0)
      raw_pkt[`PKG_SZ-18 -: `PAYLOAD_W] = payload;
  endfunction

  function void post_randomize(); 
  pack_bits(); 
  endfunction

  function string convert2str();
    return $sformatf("to[%0d,%0d] mode=%0b payload=0x%0h egress_id=%0d",
                     target_row, target_col, mode, payload, egress_id);
  endfunction
endclass
